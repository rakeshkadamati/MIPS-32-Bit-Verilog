module RegisterFile(rw,addr1,addr2,out1,out2,addr3,data3,clk);

input rw;  	//0 is read. 1 is write
input [4:0] addr1;	//rs
input [4:0] addr2;	//rt
input [4:0] addr3;	//rd
input [31:0] data3;	//value to go into addr3, rd
output [31:0] out1;	//output of read
output [31:0] out2;	//output of read


input clk;

reg [31:0] regmem [31:0]; //32x32bit array of registers

initial begin
	  regmem[0] = 32'b00000000000000000000000000000010; //2
	  regmem[1] = 32'b00000000000000000000000000000001; //1
        regmem[2] = 32'b00000000000000000000000000001000; //8
        regmem[3] = 32'b00000000000000000000000000000110; //6
        regmem[4] = 32'b00000000000000000000000001000000; //64
        regmem[5] = 32'b00000000000000000000000000100000; //32
        regmem[6] = 32'b00000000000000000000000000010000; //16
        regmem[7] = 32'b00000000000000000000000000000111; //7
        regmem[8] = 32'b00000000000000000000000000000101;  //5
        regmem[9] = 32'b00000000000000000000000000100011;  //35
        regmem[10] = 32'b00000000000000000000000000001001; //9
        regmem[11] = 32'b00000000000000000000000000001110; //14
        regmem[12] = 32'b00000000000000000000000000010010; //18
        regmem[13] = 32'b00000000000000000000000000011100; //28
        regmem[14] = 32'b00000000000000000000000000011101; //29
        regmem[15] = 32'b00000000000000000000000000001111;  //15
        regmem[16] = 32'b00000000000000000000000000001011;  //11
        regmem[17] = 32'b00000000000000000000000000010000; //16
        regmem[18] = 32'b00000000000000000000000000000001; //1
        regmem[19] = 32'b00000000000000000000000000000010; //2
        regmem[20] = 32'b00000000000000000000000000011111; //31
        regmem[21] = 32'b00000000000000000000000000010000; //16
        regmem[22] = 32'b00000000000000000000000000010001; //17
        regmem[23] = 32'b00000000000000000000000000010010; //18
        regmem[24] = 32'b00000000000000000000000000000111; //7
        regmem[25] = 32'b00000000000000000000000000111111; //63
        regmem[26] = 32'b00000000000000000000000010000000; //128
        regmem[27] = 32'b00000000000000000000000010000011; //131
        regmem[28] = 32'b00000000000000000000000000001001; //9
        regmem[29] = 32'b00000000000000000000000011000000; //192
        regmem[30] = 32'b00000000000000000000000000000111; //7
        regmem[31] = 32'b00000000000000000000000000000100; //4

	end

		assign out1 = regmem[addr1];
		assign out2 = regmem[addr2];

	//always@(rw)
	always@ (negedge clk)
	begin
		if(rw==1'b1) //if write, store data3 into addr3
		begin
		 regmem[addr3] = data3;
		end
	end

endmodule



